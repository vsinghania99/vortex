// Copyright © 2019-2023
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

interface VX_tcu_to_lsu_if ();

    wire                                valid;
    wire                                ready;
    wire [`XLEN-1:0]                    addr;   //global address in memory
    wire                                load;


    //tensor core
    modport master (
        output                          ready,
        input                           valid,
        output [`XLEN-1:0]              addr,
        output                          load;
    );

    //LSU
    modport slave (
        input                          ready,
        output                         valid,
        input [`XLEN-1:0]              addr,
        input                          load;
    );

endinterface
